library verilog;
use verilog.vl_types.all;
entity HCSR04_interface_vlg_vec_tst is
end HCSR04_interface_vlg_vec_tst;
