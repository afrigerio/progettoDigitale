library verilog;
use verilog.vl_types.all;
entity RS232_vlg_vec_tst is
end RS232_vlg_vec_tst;
