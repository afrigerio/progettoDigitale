library verilog;
use verilog.vl_types.all;
entity progetto_vlg_vec_tst is
end progetto_vlg_vec_tst;
